`timescale 1ns / 100ps

module ALU(A,B,OP,C,Cout);

	input [15:0]A;
	input [15:0]B;
	input [3:0]OP;
	output [15:0]C;
	output Cout;

	wire signed [15:0]A; 
	wire signed [15:0]B;
	wire [3:0]OP;
	reg signed [15:0]C;
	reg Cout;

	// Arithmetic
	`define	OP_ADD	4'b0000
	`define	OP_SUB	4'b0001
	// Bitwise Boolean operation
	`define	OP_AND	4'b0010
	`define	OP_OR 	4'b0011
	`define	OP_NAND	4'b0100
	`define	OP_NOR	4'b0101
	`define	OP_XOR	4'b0110
	`define	OP_XNOR	4'b0111
	// Logic
	`define	OP_ID	4'b1000
	`define	OP_NOT  4'b1001
	// Shift
	`define	OP_LRS	4'b1010
	`define	OP_ARS	4'b1011
	`define	OP_RR	4'b1100
	`define	OP_LLS	4'b1101
	`define	OP_ALS	4'b1110
	`define	OP_RL	4'b1111

	initial begin
    end

    always @(*) begin
        case (OP)
			`OP_ADD: begin
				C=A+B;
				// Overflow happens when the sign of the two operands are the same, 
				// and the sign of the output is different from the operands.
				if (A[15] ^ B[15] == 0)
					if (A[15] ^ C[15] == 1)
						Cout = 1;
					else
						Cout=0;
				else
					Cout=0;
			end

			`OP_SUB: begin
				C=A-B;
				// Overflow happens when the sign of the two operands are different, 
				// and the sign of the output is different from the first operand.
				if (A[15] ^ B[15] == 1)
					if (A[15] ^ C[15] == 1)
						Cout = 1;
					else
						Cout=0;
				else
					Cout=0;
			end

			`OP_AND: begin
				C = A&B;
				Cout = 0;
			end

			`OP_OR: begin
				C = A|B;
				Cout = 0;
			end

			`OP_NAND: begin
				C = ~(A&B);
				Cout = 0;
			end

			`OP_NOR: begin
				C = ~(A|B);
				Cout = 0;
			end

			`OP_XOR: begin
				C = A^B;
				Cout = 0;
			end

			`OP_XNOR: begin
				C = ~(A^B);
				Cout = 0;
			end

			`OP_ID: begin
				C = A;
				Cout = 0;
			end

			`OP_NOT: begin
				C = ~A;
				Cout = 0;
			end

			`OP_LRS: begin
				C = A >> 1;
				Cout = 0;
			end

			`OP_ARS: begin
				C = A >>> 1;
				Cout = 0;
			end

			`OP_RR: begin
				C = {A[0], A[15:1]};
				Cout = 0;
			end

			`OP_LLS: begin
				C = A << 1;
				Cout = 0;
			end

			`OP_ALS: begin
				C = A <<< 1;
				Cout = 0;
			end

			`OP_RL: begin
				C = {A[14:0], A[15]};
				Cout = 0;
			end

			default: begin
				C=0;
			end
		endcase
    end
	
endmodule
